library verilog;
use verilog.vl_types.all;
entity seqdec_58_t is
    generic(
        t_in_0          : integer := 26;
        t_in_1          : integer := 109896
    );
end seqdec_58_t;
