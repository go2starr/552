library verilog;
use verilog.vl_types.all;
entity quadmux4_1_t is
end quadmux4_1_t;
