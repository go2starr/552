library verilog;
use verilog.vl_types.all;
entity add4_t is
end add4_t;
