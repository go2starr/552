module detect_58_next_t();
   initial begin
      $display("Hello, world!\n");
   end
endmodule // detect_58_next_t

         

