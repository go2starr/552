library verilog;
use verilog.vl_types.all;
entity seqdec_58 is
    port(
        ina             : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        \Out\           : out    vl_logic
    );
end seqdec_58;
