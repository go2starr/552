library verilog;
use verilog.vl_types.all;
entity nor2 is
    port(
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        \out\           : out    vl_logic
    );
end nor2;
