library verilog;
use verilog.vl_types.all;
entity mux2_1_t is
end mux2_1_t;
