library verilog;
use verilog.vl_types.all;
entity detect_58_next_t is
end detect_58_next_t;
