library verilog;
use verilog.vl_types.all;
entity detect_58 is
    port(
        \in\            : in     vl_logic;
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        \out\           : out    vl_logic
    );
end detect_58;
