library verilog;
use verilog.vl_types.all;
entity fa_t is
end fa_t;
