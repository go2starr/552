library verilog;
use verilog.vl_types.all;
entity shift16_t is
end shift16_t;
