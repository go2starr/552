module detect_58_t();
   reg in, rst;

   
   
