library verilog;
use verilog.vl_types.all;
entity mux_quad4_1_t is
end mux_quad4_1_t;
