library verilog;
use verilog.vl_types.all;
entity mux4_1_t is
end mux4_1_t;
